`define DIV 2'b00
`define DIVW 2'b01
`define DIVU 2'b10
`define DIVWU 2'b11

