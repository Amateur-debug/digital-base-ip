`define UNSIGNED_X_UNSIGNED 2'b00
`define SIGNED_X_UNSIGNED 2'b01
`define SIGNED_X_SIGNED 2'b10