`timescale  1ns/1ns
module  tb_icache();

//********************************************************************//
//****************** Parameter and Internal Signal *******************//
//********************************************************************//
//parameter define
localparam RUN_TIME = 10000;

//wire  define

//reg   define

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

//initialize clock
initial begin
    clock   = 1'b0;
end
always  #10 clock = ~clock;

//initialize motivation
initial begin
	
end

always begin
    #100;
    if ($time >= RUN_TIME) begin
        $finish ;
    end
end
//********************************************************************//
//**************************** Instantiate ***************************//
//********************************************************************//

endmodule
